//Just for testing branch commits



module test();

endmodule

//some more comments for diff checking
