module test;

//just to test the git commands

endmodule